

interface adder_interface(input logic clock);

  logic reset;

  logic [7:0] input_1, input_2;
  logic [15:0] output_3;

endinterface: adder_interface
